`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Furusawa lab.
// Engineer: Ruofan He
// 
// Create Date: 2021/10/21 18:03:08
// Design Name: 
// Module Name: PNR_register
// Project Name: redpitaya_PNR
// Target Devices:
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PNR_register(
   // signals
   input  wire            clk_i           ,  //!< processing clock
   input  wire            rstn_i          ,  //!< processing reset - active low

   //led test
   output reg [8-1:0]    led_o           ,
   // system bus
   input  wire [ 32-1: 0] sys_addr        ,  //!< bus address
   input  wire [ 32-1: 0] sys_wdata       ,  //!< bus write data
   input  wire            sys_wen         ,  //!< bus write enable
   input  wire            sys_ren         ,  //!< bus read enable
   output reg [ 32-1: 0] sys_rdata       ,  //!< bus read data
   output reg            sys_err         ,  //!< bus error indicator
   output reg            sys_ack         ,  //!< bus acknowledge signal
   //ADC_threshold for photon number resolving
   output reg [ 14-1: 0] adc_photon_threshold_1,
   output reg [ 14-1: 0] adc_photon_threshold_2,
   output reg [ 14-1: 0] adc_photon_threshold_3,
   output reg [ 14-1: 0] adc_photon_threshold_4,
   output reg [ 14-1: 0] adc_photon_threshold_5,
   output reg [ 14-1: 0] adc_photon_threshold_6,
   output reg [ 14-1: 0] adc_photon_threshold_7
    );

//---------------------------------------------------------------------------------
//
//  System bus connection

always @(posedge clk_i) begin
   if (rstn_i == 1'b0) begin
      led_o    <= 8'h0 ;
      adc_photon_threshold_1  <= 14'b0;
      adc_photon_threshold_2  <= 14'b0;
      adc_photon_threshold_3  <= 14'b0;
      adc_photon_threshold_4  <= 14'b0;
      adc_photon_threshold_5  <= 14'b0;
      adc_photon_threshold_6  <= 14'b0;
      adc_photon_threshold_7  <= 14'b0;

   end
   else begin
      if (sys_wen) begin
         if (sys_addr[20-1:0]==20'h00)    led_o  <= sys_wdata[8-1:0] ;
         if (sys_addr[20-1:0]==20'h04)    adc_photon_threshold_1  <= sys_wdata[14-1:0] ;
         if (sys_addr[20-1:0]==20'h08)    adc_photon_threshold_2  <= sys_wdata[14-1:0] ;
         if (sys_addr[20-1:0]==20'h0C)    adc_photon_threshold_3  <= sys_wdata[14-1:0] ;
         if (sys_addr[20-1:0]==20'h10)    adc_photon_threshold_4  <= sys_wdata[14-1:0] ;
         if (sys_addr[20-1:0]==20'h14)    adc_photon_threshold_5  <= sys_wdata[14-1:0] ;
         if (sys_addr[20-1:0]==20'h18)    adc_photon_threshold_6  <= sys_wdata[14-1:0] ;
         if (sys_addr[20-1:0]==20'h1C)    adc_photon_threshold_7  <= sys_wdata[14-1:0] ;
      end
   end
end

wire sys_en;
assign sys_en = sys_wen | sys_ren;

always @(posedge clk_i)
if (rstn_i == 1'b0) begin
   sys_err <= 1'b0 ;
   sys_ack <= 1'b0 ;
end else begin
   sys_err <= 1'b0 ;

   casez (sys_addr[20-1:0])
      20'h00  : begin sys_ack <= sys_en;         sys_rdata <= {{32- 8{1'b00}}, led_o                 }              ; end
      20'h04  : begin sys_ack <= sys_en;         sys_rdata <= {{32-14{1'b04}}, adc_photon_threshold_1}              ; end
      20'h08  : begin sys_ack <= sys_en;         sys_rdata <= {{32-14{1'b08}}, adc_photon_threshold_2}              ; end
      20'h0C  : begin sys_ack <= sys_en;         sys_rdata <= {{32-14{1'b0C}}, adc_photon_threshold_3}              ; end
      20'h10  : begin sys_ack <= sys_en;         sys_rdata <= {{32-14{1'b10}}, adc_photon_threshold_4}              ; end
      20'h14  : begin sys_ack <= sys_en;         sys_rdata <= {{32-14{1'b14}}, adc_photon_threshold_5}              ; end
      20'h18  : begin sys_ack <= sys_en;         sys_rdata <= {{32-14{1'b18}}, adc_photon_threshold_6}              ; end
      20'h1C  : begin sys_ack <= sys_en;         sys_rdata <= {{32-14{1'b1C}}, adc_photon_threshold_7}              ; end
      default : begin sys_ack <= sys_en;         sys_rdata <=  32'h0                                                ; end
   endcase
end

endmodule

